/*
* Piggy Bank
* Adds credit for penny(1), nickel(5), dime(10), and quarter(25)
* Subtracts credit for apple(75), banana(20), carrot(30), and date(40)
* Max credit is $2.55, displayed in hex
* Resets asynchronously
*/

module piggyBank (input clk, reset, penny, nickel, dime, quarter, apple, banana, carrot, date, output [7:0] credit);
  input clk, reset, penny, nickel, dime, quarter, apple, banana, carrot, date;
  output [7:0] credit;
  
  always @ (posedge clk or reset)
  
  begin
  
  
  
  
  
  
  end
endmodule
