module coinSensor(penny,nickel,dime,quarter, clk,reset,serialIn);
  output penny, nickel, dime, quarter;
  input clk, reset, serialIn;
  
  





endmodule
